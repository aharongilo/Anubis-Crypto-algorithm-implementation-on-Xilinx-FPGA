
module mult_rom8
(
	input [7:0]data_in,
	output reg [7:0] data_out
);
always@(data_in)
    case (data_in)  
				0 : data_out <=8'h0;
		1 : data_out <=8'h8;
		2 : data_out <=8'h10;
		3 : data_out <=8'h18;
		4 : data_out <=8'h20;
		5 : data_out <=8'h28;
		6 : data_out <=8'h30;
		7 : data_out <=8'h38;
		8 : data_out <=8'h40;
		9 : data_out <=8'h48;
		10 : data_out <=8'h50;
		11 : data_out <=8'h58;
		12 : data_out <=8'h60;
		13 : data_out <=8'h68;
		14 : data_out <=8'h70;
		15 : data_out <=8'h78;
		16 : data_out <=8'h80;
		17 : data_out <=8'h88;
		18 : data_out <=8'h90;
		19 : data_out <=8'h98;
		20 : data_out <=8'ha0;
		21 : data_out <=8'ha8;
		22 : data_out <=8'hb0;
		23 : data_out <=8'hb8;
		24 : data_out <=8'hc0;
		25 : data_out <=8'hc8;
		26 : data_out <=8'hd0;
		27 : data_out <=8'hd8;
		28 : data_out <=8'he0;
		29 : data_out <=8'he8;
		30 : data_out <=8'hf0;
		31 : data_out <=8'hf8;
		32 : data_out <=8'h1d;
		33 : data_out <=8'h15;
		34 : data_out <=8'hd;
		35 : data_out <=8'h5;
		36 : data_out <=8'h3d;
		37 : data_out <=8'h35;
		38 : data_out <=8'h2d;
		39 : data_out <=8'h25;
		40 : data_out <=8'h5d;
		41 : data_out <=8'h55;
		42 : data_out <=8'h4d;
		43 : data_out <=8'h45;
		44 : data_out <=8'h7d;
		45 : data_out <=8'h75;
		46 : data_out <=8'h6d;
		47 : data_out <=8'h65;
		48 : data_out <=8'h9d;
		49 : data_out <=8'h95;
		50 : data_out <=8'h8d;
		51 : data_out <=8'h85;
		52 : data_out <=8'hbd;
		53 : data_out <=8'hb5;
		54 : data_out <=8'had;
		55 : data_out <=8'ha5;
		56 : data_out <=8'hdd;
		57 : data_out <=8'hd5;
		58 : data_out <=8'hcd;
		59 : data_out <=8'hc5;
		60 : data_out <=8'hfd;
		61 : data_out <=8'hf5;
		62 : data_out <=8'hed;
		63 : data_out <=8'he5;
		64 : data_out <=8'h3a;
		65 : data_out <=8'h32;
		66 : data_out <=8'h2a;
		67 : data_out <=8'h22;
		68 : data_out <=8'h1a;
		69 : data_out <=8'h12;
		70 : data_out <=8'ha;
		71 : data_out <=8'h2;
		72 : data_out <=8'h7a;
		73 : data_out <=8'h72;
		74 : data_out <=8'h6a;
		75 : data_out <=8'h62;
		76 : data_out <=8'h5a;
		77 : data_out <=8'h52;
		78 : data_out <=8'h4a;
		79 : data_out <=8'h42;
		80 : data_out <=8'hba;
		81 : data_out <=8'hb2;
		82 : data_out <=8'haa;
		83 : data_out <=8'ha2;
		84 : data_out <=8'h9a;
		85 : data_out <=8'h92;
		86 : data_out <=8'h8a;
		87 : data_out <=8'h82;
		88 : data_out <=8'hfa;
		89 : data_out <=8'hf2;
		90 : data_out <=8'hea;
		91 : data_out <=8'he2;
		92 : data_out <=8'hda;
		93 : data_out <=8'hd2;
		94 : data_out <=8'hca;
		95 : data_out <=8'hc2;
		96 : data_out <=8'h27;
		97 : data_out <=8'h2f;
		98 : data_out <=8'h37;
		99 : data_out <=8'h3f;
		100 : data_out <=8'h7;
		101 : data_out <=8'hf;
		102 : data_out <=8'h17;
		103 : data_out <=8'h1f;
		104 : data_out <=8'h67;
		105 : data_out <=8'h6f;
		106 : data_out <=8'h77;
		107 : data_out <=8'h7f;
		108 : data_out <=8'h47;
		109 : data_out <=8'h4f;
		110 : data_out <=8'h57;
		111 : data_out <=8'h5f;
		112 : data_out <=8'ha7;
		113 : data_out <=8'haf;
		114 : data_out <=8'hb7;
		115 : data_out <=8'hbf;
		116 : data_out <=8'h87;
		117 : data_out <=8'h8f;
		118 : data_out <=8'h97;
		119 : data_out <=8'h9f;
		120 : data_out <=8'he7;
		121 : data_out <=8'hef;
		122 : data_out <=8'hf7;
		123 : data_out <=8'hff;
		124 : data_out <=8'hc7;
		125 : data_out <=8'hcf;
		126 : data_out <=8'hd7;
		127 : data_out <=8'hdf;
		128 : data_out <=8'h74;
		129 : data_out <=8'h7c;
		130 : data_out <=8'h64;
		131 : data_out <=8'h6c;
		132 : data_out <=8'h54;
		133 : data_out <=8'h5c;
		134 : data_out <=8'h44;
		135 : data_out <=8'h4c;
		136 : data_out <=8'h34;
		137 : data_out <=8'h3c;
		138 : data_out <=8'h24;
		139 : data_out <=8'h2c;
		140 : data_out <=8'h14;
		141 : data_out <=8'h1c;
		142 : data_out <=8'h4;
		143 : data_out <=8'hc;
		144 : data_out <=8'hf4;
		145 : data_out <=8'hfc;
		146 : data_out <=8'he4;
		147 : data_out <=8'hec;
		148 : data_out <=8'hd4;
		149 : data_out <=8'hdc;
		150 : data_out <=8'hc4;
		151 : data_out <=8'hcc;
		152 : data_out <=8'hb4;
		153 : data_out <=8'hbc;
		154 : data_out <=8'ha4;
		155 : data_out <=8'hac;
		156 : data_out <=8'h94;
		157 : data_out <=8'h9c;
		158 : data_out <=8'h84;
		159 : data_out <=8'h8c;
		160 : data_out <=8'h69;
		161 : data_out <=8'h61;
		162 : data_out <=8'h79;
		163 : data_out <=8'h71;
		164 : data_out <=8'h49;
		165 : data_out <=8'h41;
		166 : data_out <=8'h59;
		167 : data_out <=8'h51;
		168 : data_out <=8'h29;
		169 : data_out <=8'h21;
		170 : data_out <=8'h39;
		171 : data_out <=8'h31;
		172 : data_out <=8'h9;
		173 : data_out <=8'h1;
		174 : data_out <=8'h19;
		175 : data_out <=8'h11;
		176 : data_out <=8'he9;
		177 : data_out <=8'he1;
		178 : data_out <=8'hf9;
		179 : data_out <=8'hf1;
		180 : data_out <=8'hc9;
		181 : data_out <=8'hc1;
		182 : data_out <=8'hd9;
		183 : data_out <=8'hd1;
		184 : data_out <=8'ha9;
		185 : data_out <=8'ha1;
		186 : data_out <=8'hb9;
		187 : data_out <=8'hb1;
		188 : data_out <=8'h89;
		189 : data_out <=8'h81;
		190 : data_out <=8'h99;
		191 : data_out <=8'h91;
		192 : data_out <=8'h4e;
		193 : data_out <=8'h46;
		194 : data_out <=8'h5e;
		195 : data_out <=8'h56;
		196 : data_out <=8'h6e;
		197 : data_out <=8'h66;
		198 : data_out <=8'h7e;
		199 : data_out <=8'h76;
		200 : data_out <=8'he;
		201 : data_out <=8'h6;
		202 : data_out <=8'h1e;
		203 : data_out <=8'h16;
		204 : data_out <=8'h2e;
		205 : data_out <=8'h26;
		206 : data_out <=8'h3e;
		207 : data_out <=8'h36;
		208 : data_out <=8'hce;
		209 : data_out <=8'hc6;
		210 : data_out <=8'hde;
		211 : data_out <=8'hd6;
		212 : data_out <=8'hee;
		213 : data_out <=8'he6;
		214 : data_out <=8'hfe;
		215 : data_out <=8'hf6;
		216 : data_out <=8'h8e;
		217 : data_out <=8'h86;
		218 : data_out <=8'h9e;
		219 : data_out <=8'h96;
		220 : data_out <=8'hae;
		221 : data_out <=8'ha6;
		222 : data_out <=8'hbe;
		223 : data_out <=8'hb6;
		224 : data_out <=8'h53;
		225 : data_out <=8'h5b;
		226 : data_out <=8'h43;
		227 : data_out <=8'h4b;
		228 : data_out <=8'h73;
		229 : data_out <=8'h7b;
		230 : data_out <=8'h63;
		231 : data_out <=8'h6b;
		232 : data_out <=8'h13;
		233 : data_out <=8'h1b;
		234 : data_out <=8'h3;
		235 : data_out <=8'hb;
		236 : data_out <=8'h33;
		237 : data_out <=8'h3b;
		238 : data_out <=8'h23;
		239 : data_out <=8'h2b;
		240 : data_out <=8'hd3;
		241 : data_out <=8'hdb;
		242 : data_out <=8'hc3;
		243 : data_out <=8'hcb;
		244 : data_out <=8'hf3;
		245 : data_out <=8'hfb;
		246 : data_out <=8'he3;
		247 : data_out <=8'heb;
		248 : data_out <=8'h93;
		249 : data_out <=8'h9b;
		250 : data_out <=8'h83;
		251 : data_out <=8'h8b;
		252 : data_out <=8'hb3;
		253 : data_out <=8'hbb;
		254 : data_out <=8'ha3;
		255 : data_out <=8'hab;

		default: data_out<= 8'h0;
    endcase

endmodule
