
module mult_rom2
(
	input [7:0]data_in,
	output reg [7:0] data_out
);
always@(data_in)
    case (data_in)  
		0 : data_out <=8'h0;
		1 : data_out <=8'h2;
		2 : data_out <=8'h4;
		3 : data_out <=8'h6;
		4 : data_out <=8'h8;
		5 : data_out <=8'ha;
		6 : data_out <=8'hc;
		7 : data_out <=8'he;
		8 : data_out <=8'h10;
		9 : data_out <=8'h12;
		10 : data_out <=8'h14;
		11 : data_out <=8'h16;
		12 : data_out <=8'h18;
		13 : data_out <=8'h1a;
		14 : data_out <=8'h1c;
		15 : data_out <=8'h1e;
		16 : data_out <=8'h20;
		17 : data_out <=8'h22;
		18 : data_out <=8'h24;
		19 : data_out <=8'h26;
		20 : data_out <=8'h28;
		21 : data_out <=8'h2a;
		22 : data_out <=8'h2c;
		23 : data_out <=8'h2e;
		24 : data_out <=8'h30;
		25 : data_out <=8'h32;
		26 : data_out <=8'h34;
		27 : data_out <=8'h36;
		28 : data_out <=8'h38;
		29 : data_out <=8'h3a;
		30 : data_out <=8'h3c;
		31 : data_out <=8'h3e;
		32 : data_out <=8'h40;
		33 : data_out <=8'h42;
		34 : data_out <=8'h44;
		35 : data_out <=8'h46;
		36 : data_out <=8'h48;
		37 : data_out <=8'h4a;
		38 : data_out <=8'h4c;
		39 : data_out <=8'h4e;
		40 : data_out <=8'h50;
		41 : data_out <=8'h52;
		42 : data_out <=8'h54;
		43 : data_out <=8'h56;
		44 : data_out <=8'h58;
		45 : data_out <=8'h5a;
		46 : data_out <=8'h5c;
		47 : data_out <=8'h5e;
		48 : data_out <=8'h60;
		49 : data_out <=8'h62;
		50 : data_out <=8'h64;
		51 : data_out <=8'h66;
		52 : data_out <=8'h68;
		53 : data_out <=8'h6a;
		54 : data_out <=8'h6c;
		55 : data_out <=8'h6e;
		56 : data_out <=8'h70;
		57 : data_out <=8'h72;
		58 : data_out <=8'h74;
		59 : data_out <=8'h76;
		60 : data_out <=8'h78;
		61 : data_out <=8'h7a;
		62 : data_out <=8'h7c;
		63 : data_out <=8'h7e;
		64 : data_out <=8'h80;
		65 : data_out <=8'h82;
		66 : data_out <=8'h84;
		67 : data_out <=8'h86;
		68 : data_out <=8'h88;
		69 : data_out <=8'h8a;
		70 : data_out <=8'h8c;
		71 : data_out <=8'h8e;
		72 : data_out <=8'h90;
		73 : data_out <=8'h92;
		74 : data_out <=8'h94;
		75 : data_out <=8'h96;
		76 : data_out <=8'h98;
		77 : data_out <=8'h9a;
		78 : data_out <=8'h9c;
		79 : data_out <=8'h9e;
		80 : data_out <=8'ha0;
		81 : data_out <=8'ha2;
		82 : data_out <=8'ha4;
		83 : data_out <=8'ha6;
		84 : data_out <=8'ha8;
		85 : data_out <=8'haa;
		86 : data_out <=8'hac;
		87 : data_out <=8'hae;
		88 : data_out <=8'hb0;
		89 : data_out <=8'hb2;
		90 : data_out <=8'hb4;
		91 : data_out <=8'hb6;
		92 : data_out <=8'hb8;
		93 : data_out <=8'hba;
		94 : data_out <=8'hbc;
		95 : data_out <=8'hbe;
		96 : data_out <=8'hc0;
		97 : data_out <=8'hc2;
		98 : data_out <=8'hc4;
		99 : data_out <=8'hc6;
		100 : data_out <=8'hc8;
		101 : data_out <=8'hca;
		102 : data_out <=8'hcc;
		103 : data_out <=8'hce;
		104 : data_out <=8'hd0;
		105 : data_out <=8'hd2;
		106 : data_out <=8'hd4;
		107 : data_out <=8'hd6;
		108 : data_out <=8'hd8;
		109 : data_out <=8'hda;
		110 : data_out <=8'hdc;
		111 : data_out <=8'hde;
		112 : data_out <=8'he0;
		113 : data_out <=8'he2;
		114 : data_out <=8'he4;
		115 : data_out <=8'he6;
		116 : data_out <=8'he8;
		117 : data_out <=8'hea;
		118 : data_out <=8'hec;
		119 : data_out <=8'hee;
		120 : data_out <=8'hf0;
		121 : data_out <=8'hf2;
		122 : data_out <=8'hf4;
		123 : data_out <=8'hf6;
		124 : data_out <=8'hf8;
		125 : data_out <=8'hfa;
		126 : data_out <=8'hfc;
		127 : data_out <=8'hfe;
		128 : data_out <=8'h1d;
		129 : data_out <=8'h1f;
		130 : data_out <=8'h19;
		131 : data_out <=8'h1b;
		132 : data_out <=8'h15;
		133 : data_out <=8'h17;
		134 : data_out <=8'h11;
		135 : data_out <=8'h13;
		136 : data_out <=8'hd;
		137 : data_out <=8'hf;
		138 : data_out <=8'h9;
		139 : data_out <=8'hb;
		140 : data_out <=8'h5;
		141 : data_out <=8'h7;
		142 : data_out <=8'h1;
		143 : data_out <=8'h3;
		144 : data_out <=8'h3d;
		145 : data_out <=8'h3f;
		146 : data_out <=8'h39;
		147 : data_out <=8'h3b;
		148 : data_out <=8'h35;
		149 : data_out <=8'h37;
		150 : data_out <=8'h31;
		151 : data_out <=8'h33;
		152 : data_out <=8'h2d;
		153 : data_out <=8'h2f;
		154 : data_out <=8'h29;
		155 : data_out <=8'h2b;
		156 : data_out <=8'h25;
		157 : data_out <=8'h27;
		158 : data_out <=8'h21;
		159 : data_out <=8'h23;
		160 : data_out <=8'h5d;
		161 : data_out <=8'h5f;
		162 : data_out <=8'h59;
		163 : data_out <=8'h5b;
		164 : data_out <=8'h55;
		165 : data_out <=8'h57;
		166 : data_out <=8'h51;
		167 : data_out <=8'h53;
		168 : data_out <=8'h4d;
		169 : data_out <=8'h4f;
		170 : data_out <=8'h49;
		171 : data_out <=8'h4b;
		172 : data_out <=8'h45;
		173 : data_out <=8'h47;
		174 : data_out <=8'h41;
		175 : data_out <=8'h43;
		176 : data_out <=8'h7d;
		177 : data_out <=8'h7f;
		178 : data_out <=8'h79;
		179 : data_out <=8'h7b;
		180 : data_out <=8'h75;
		181 : data_out <=8'h77;
		182 : data_out <=8'h71;
		183 : data_out <=8'h73;
		184 : data_out <=8'h6d;
		185 : data_out <=8'h6f;
		186 : data_out <=8'h69;
		187 : data_out <=8'h6b;
		188 : data_out <=8'h65;
		189 : data_out <=8'h67;
		190 : data_out <=8'h61;
		191 : data_out <=8'h63;
		192 : data_out <=8'h9d;
		193 : data_out <=8'h9f;
		194 : data_out <=8'h99;
		195 : data_out <=8'h9b;
		196 : data_out <=8'h95;
		197 : data_out <=8'h97;
		198 : data_out <=8'h91;
		199 : data_out <=8'h93;
		200 : data_out <=8'h8d;
		201 : data_out <=8'h8f;
		202 : data_out <=8'h89;
		203 : data_out <=8'h8b;
		204 : data_out <=8'h85;
		205 : data_out <=8'h87;
		206 : data_out <=8'h81;
		207 : data_out <=8'h83;
		208 : data_out <=8'hbd;
		209 : data_out <=8'hbf;
		210 : data_out <=8'hb9;
		211 : data_out <=8'hbb;
		212 : data_out <=8'hb5;
		213 : data_out <=8'hb7;
		214 : data_out <=8'hb1;
		215 : data_out <=8'hb3;
		216 : data_out <=8'had;
		217 : data_out <=8'haf;
		218 : data_out <=8'ha9;
		219 : data_out <=8'hab;
		220 : data_out <=8'ha5;
		221 : data_out <=8'ha7;
		222 : data_out <=8'ha1;
		223 : data_out <=8'ha3;
		224 : data_out <=8'hdd;
		225 : data_out <=8'hdf;
		226 : data_out <=8'hd9;
		227 : data_out <=8'hdb;
		228 : data_out <=8'hd5;
		229 : data_out <=8'hd7;
		230 : data_out <=8'hd1;
		231 : data_out <=8'hd3;
		232 : data_out <=8'hcd;
		233 : data_out <=8'hcf;
		234 : data_out <=8'hc9;
		235 : data_out <=8'hcb;
		236 : data_out <=8'hc5;
		237 : data_out <=8'hc7;
		238 : data_out <=8'hc1;
		239 : data_out <=8'hc3;
		240 : data_out <=8'hfd;
		241 : data_out <=8'hff;
		242 : data_out <=8'hf9;
		243 : data_out <=8'hfb;
		244 : data_out <=8'hf5;
		245 : data_out <=8'hf7;
		246 : data_out <=8'hf1;
		247 : data_out <=8'hf3;
		248 : data_out <=8'hed;
		249 : data_out <=8'hef;
		250 : data_out <=8'he9;
		251 : data_out <=8'heb;
		252 : data_out <=8'he5;
		253 : data_out <=8'he7;
		254 : data_out <=8'he1;
		255 : data_out <=8'he3;
		default: data_out<= 8'h0;
    endcase

endmodule
