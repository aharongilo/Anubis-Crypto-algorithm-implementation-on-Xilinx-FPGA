
module mult_rom4
(
	input [7:0]data_in,
	output reg [7:0] data_out
);
always@(data_in)
    case (data_in)  
		0 : data_out <=8'h0;
		1 : data_out <=8'h4;
		2 : data_out <=8'h8;
		3 : data_out <=8'hc;
		4 : data_out <=8'h10;
		5 : data_out <=8'h14;
		6 : data_out <=8'h18;
		7 : data_out <=8'h1c;
		8 : data_out <=8'h20;
		9 : data_out <=8'h24;
		10 : data_out <=8'h28;
		11 : data_out <=8'h2c;
		12 : data_out <=8'h30;
		13 : data_out <=8'h34;
		14 : data_out <=8'h38;
		15 : data_out <=8'h3c;
		16 : data_out <=8'h40;
		17 : data_out <=8'h44;
		18 : data_out <=8'h48;
		19 : data_out <=8'h4c;
		20 : data_out <=8'h50;
		21 : data_out <=8'h54;
		22 : data_out <=8'h58;
		23 : data_out <=8'h5c;
		24 : data_out <=8'h60;
		25 : data_out <=8'h64;
		26 : data_out <=8'h68;
		27 : data_out <=8'h6c;
		28 : data_out <=8'h70;
		29 : data_out <=8'h74;
		30 : data_out <=8'h78;
		31 : data_out <=8'h7c;
		32 : data_out <=8'h80;
		33 : data_out <=8'h84;
		34 : data_out <=8'h88;
		35 : data_out <=8'h8c;
		36 : data_out <=8'h90;
		37 : data_out <=8'h94;
		38 : data_out <=8'h98;
		39 : data_out <=8'h9c;
		40 : data_out <=8'ha0;
		41 : data_out <=8'ha4;
		42 : data_out <=8'ha8;
		43 : data_out <=8'hac;
		44 : data_out <=8'hb0;
		45 : data_out <=8'hb4;
		46 : data_out <=8'hb8;
		47 : data_out <=8'hbc;
		48 : data_out <=8'hc0;
		49 : data_out <=8'hc4;
		50 : data_out <=8'hc8;
		51 : data_out <=8'hcc;
		52 : data_out <=8'hd0;
		53 : data_out <=8'hd4;
		54 : data_out <=8'hd8;
		55 : data_out <=8'hdc;
		56 : data_out <=8'he0;
		57 : data_out <=8'he4;
		58 : data_out <=8'he8;
		59 : data_out <=8'hec;
		60 : data_out <=8'hf0;
		61 : data_out <=8'hf4;
		62 : data_out <=8'hf8;
		63 : data_out <=8'hfc;
		64 : data_out <=8'h1d;
		65 : data_out <=8'h19;
		66 : data_out <=8'h15;
		67 : data_out <=8'h11;
		68 : data_out <=8'hd;
		69 : data_out <=8'h9;
		70 : data_out <=8'h5;
		71 : data_out <=8'h1;
		72 : data_out <=8'h3d;
		73 : data_out <=8'h39;
		74 : data_out <=8'h35;
		75 : data_out <=8'h31;
		76 : data_out <=8'h2d;
		77 : data_out <=8'h29;
		78 : data_out <=8'h25;
		79 : data_out <=8'h21;
		80 : data_out <=8'h5d;
		81 : data_out <=8'h59;
		82 : data_out <=8'h55;
		83 : data_out <=8'h51;
		84 : data_out <=8'h4d;
		85 : data_out <=8'h49;
		86 : data_out <=8'h45;
		87 : data_out <=8'h41;
		88 : data_out <=8'h7d;
		89 : data_out <=8'h79;
		90 : data_out <=8'h75;
		91 : data_out <=8'h71;
		92 : data_out <=8'h6d;
		93 : data_out <=8'h69;
		94 : data_out <=8'h65;
		95 : data_out <=8'h61;
		96 : data_out <=8'h9d;
		97 : data_out <=8'h99;
		98 : data_out <=8'h95;
		99 : data_out <=8'h91;
		100 : data_out <=8'h8d;
		101 : data_out <=8'h89;
		102 : data_out <=8'h85;
		103 : data_out <=8'h81;
		104 : data_out <=8'hbd;
		105 : data_out <=8'hb9;
		106 : data_out <=8'hb5;
		107 : data_out <=8'hb1;
		108 : data_out <=8'had;
		109 : data_out <=8'ha9;
		110 : data_out <=8'ha5;
		111 : data_out <=8'ha1;
		112 : data_out <=8'hdd;
		113 : data_out <=8'hd9;
		114 : data_out <=8'hd5;
		115 : data_out <=8'hd1;
		116 : data_out <=8'hcd;
		117 : data_out <=8'hc9;
		118 : data_out <=8'hc5;
		119 : data_out <=8'hc1;
		120 : data_out <=8'hfd;
		121 : data_out <=8'hf9;
		122 : data_out <=8'hf5;
		123 : data_out <=8'hf1;
		124 : data_out <=8'hed;
		125 : data_out <=8'he9;
		126 : data_out <=8'he5;
		127 : data_out <=8'he1;
		128 : data_out <=8'h3a;
		129 : data_out <=8'h3e;
		130 : data_out <=8'h32;
		131 : data_out <=8'h36;
		132 : data_out <=8'h2a;
		133 : data_out <=8'h2e;
		134 : data_out <=8'h22;
		135 : data_out <=8'h26;
		136 : data_out <=8'h1a;
		137 : data_out <=8'h1e;
		138 : data_out <=8'h12;
		139 : data_out <=8'h16;
		140 : data_out <=8'ha;
		141 : data_out <=8'he;
		142 : data_out <=8'h2;
		143 : data_out <=8'h6;
		144 : data_out <=8'h7a;
		145 : data_out <=8'h7e;
		146 : data_out <=8'h72;
		147 : data_out <=8'h76;
		148 : data_out <=8'h6a;
		149 : data_out <=8'h6e;
		150 : data_out <=8'h62;
		151 : data_out <=8'h66;
		152 : data_out <=8'h5a;
		153 : data_out <=8'h5e;
		154 : data_out <=8'h52;
		155 : data_out <=8'h56;
		156 : data_out <=8'h4a;
		157 : data_out <=8'h4e;
		158 : data_out <=8'h42;
		159 : data_out <=8'h46;
		160 : data_out <=8'hba;
		161 : data_out <=8'hbe;
		162 : data_out <=8'hb2;
		163 : data_out <=8'hb6;
		164 : data_out <=8'haa;
		165 : data_out <=8'hae;
		166 : data_out <=8'ha2;
		167 : data_out <=8'ha6;
		168 : data_out <=8'h9a;
		169 : data_out <=8'h9e;
		170 : data_out <=8'h92;
		171 : data_out <=8'h96;
		172 : data_out <=8'h8a;
		173 : data_out <=8'h8e;
		174 : data_out <=8'h82;
		175 : data_out <=8'h86;
		176 : data_out <=8'hfa;
		177 : data_out <=8'hfe;
		178 : data_out <=8'hf2;
		179 : data_out <=8'hf6;
		180 : data_out <=8'hea;
		181 : data_out <=8'hee;
		182 : data_out <=8'he2;
		183 : data_out <=8'he6;
		184 : data_out <=8'hda;
		185 : data_out <=8'hde;
		186 : data_out <=8'hd2;
		187 : data_out <=8'hd6;
		188 : data_out <=8'hca;
		189 : data_out <=8'hce;
		190 : data_out <=8'hc2;
		191 : data_out <=8'hc6;
		192 : data_out <=8'h27;
		193 : data_out <=8'h23;
		194 : data_out <=8'h2f;
		195 : data_out <=8'h2b;
		196 : data_out <=8'h37;
		197 : data_out <=8'h33;
		198 : data_out <=8'h3f;
		199 : data_out <=8'h3b;
		200 : data_out <=8'h7;
		201 : data_out <=8'h3;
		202 : data_out <=8'hf;
		203 : data_out <=8'hb;
		204 : data_out <=8'h17;
		205 : data_out <=8'h13;
		206 : data_out <=8'h1f;
		207 : data_out <=8'h1b;
		208 : data_out <=8'h67;
		209 : data_out <=8'h63;
		210 : data_out <=8'h6f;
		211 : data_out <=8'h6b;
		212 : data_out <=8'h77;
		213 : data_out <=8'h73;
		214 : data_out <=8'h7f;
		215 : data_out <=8'h7b;
		216 : data_out <=8'h47;
		217 : data_out <=8'h43;
		218 : data_out <=8'h4f;
		219 : data_out <=8'h4b;
		220 : data_out <=8'h57;
		221 : data_out <=8'h53;
		222 : data_out <=8'h5f;
		223 : data_out <=8'h5b;
		224 : data_out <=8'ha7;
		225 : data_out <=8'ha3;
		226 : data_out <=8'haf;
		227 : data_out <=8'hab;
		228 : data_out <=8'hb7;
		229 : data_out <=8'hb3;
		230 : data_out <=8'hbf;
		231 : data_out <=8'hbb;
		232 : data_out <=8'h87;
		233 : data_out <=8'h83;
		234 : data_out <=8'h8f;
		235 : data_out <=8'h8b;
		236 : data_out <=8'h97;
		237 : data_out <=8'h93;
		238 : data_out <=8'h9f;
		239 : data_out <=8'h9b;
		240 : data_out <=8'he7;
		241 : data_out <=8'he3;
		242 : data_out <=8'hef;
		243 : data_out <=8'heb;
		244 : data_out <=8'hf7;
		245 : data_out <=8'hf3;
		246 : data_out <=8'hff;
		247 : data_out <=8'hfb;
		248 : data_out <=8'hc7;
		249 : data_out <=8'hc3;
		250 : data_out <=8'hcf;
		251 : data_out <=8'hcb;
		252 : data_out <=8'hd7;
		253 : data_out <=8'hd3;
		254 : data_out <=8'hdf;
		255 : data_out <=8'hdb;

		default: data_out<= 8'h0;
    endcase

endmodule
